package test_pkg;
`include "uvm_macros.svh"
import uvm_pkg::*;

`include "uvm_macros.svh"

`include "seq_item.sv"
`include "base_seq.sv"
`include "driver.sv"
`include "monitor.sv"
`include "sequencer.sv"
`include "agent.sv"
`include "scoreboaed.sv"
`include "env.sv"
`include "test.sv"

endpackage

